module microprocessor();

endmodule
