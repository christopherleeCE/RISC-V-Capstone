// This is the former memory module but renamed as the data memory
// This should function as a RAM due to its option to write to it
// A similar, read-only module has been created as the instruction memory

module data_memory
  #( 
     parameter int BIT_WIDTH,
     parameter int ENTRY_COUNT,
     parameter int ADDR_WIDTH=32 //I think this is correct for byte-addressable mem. 
     )
   (
    input  logic [ADDR_WIDTH-1:0] readAddr,
    input  logic [ADDR_WIDTH-1:0] writeAddr,
    input  logic [BIT_WIDTH-1:0] writeData,
    input  logic          writeEn,
    output logic [BIT_WIDTH-1:0] readData,
    input  logic          clk
    );

   logic [BIT_WIDTH-1:0] data_mem [ENTRY_COUNT-1:0];

   //Need this to initialize the memory
   initial begin
    $readmemh("data_memory.txt", data_mem); //load the memory
   end

   assign readData = data_mem[readAddr[ADDR_WIDTH-1:2]];

   always @(posedge clk) begin
      if( writeEn == 1'b1) begin
          data_mem[writeAddr[ADDR_WIDTH-1:2]] <= writeData ; // probably should be non-blocking
      end
   end

   
endmodule 
    