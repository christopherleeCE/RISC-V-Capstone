/*
TESTING: ADD, OR, AND

We can have a main TB for the CPU if we really need to, but I like the idea of splitting the TB for each instruction type.
In theory, each type will have a similar datapath, so in theory, each type can use a similar verification process, I'll
have to see for sure though.

I have a couple ideas for a TB but I have to figure out the implementation and see if it works. I'll be focused on these
three instructions for now; to others doing verification, please feel free to test the other instructions, thank you!



*/

module r_type_tb ();

endmodule