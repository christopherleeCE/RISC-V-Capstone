module top_register_file();

endmodule