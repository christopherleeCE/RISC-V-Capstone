module top_alu
#()
();

endmodule